module day16

pub fn task1() string {
	return "?"
}

pub fn task2() string { 
        return "?"
}

