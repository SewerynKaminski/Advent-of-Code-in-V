module day22

pub fn task1() string {
	return "1"
}

pub fn task2() string { 
        return "2"
}

